rom_sigmoid_inst : rom_sigmoid PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
