library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;  

entity network is --main entity
    port (
      clk : in std_logic;
      rst : in std_logic
      );
end entity;

architecture network_rtl of network is


begin


end architecture;